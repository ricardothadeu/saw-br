module teste_placa (
  input [3:0] entradas,
    output [3:0] saidas
);

    assign saidas = entradas;

endmodule
