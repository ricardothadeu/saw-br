module font_rom (
    input  wire [7:0] char_code,   // caractere ASCII
    input  wire [2:0] row,         // linha do caractere (0 a 7)
    output reg  [7:0] pixels       // pixels da linha (1 = ligado)
);
    always @(*) begin
        case (char_code)
            // Código ASCII das letras usadas: P R O G A M   C U N T E
            "P": case(row) 8'b11110000,8'b10001000,8'b11110000,8'b10000000,8'b10000000,8'b10000000,8'b00000000,8'b00000000; endcase
            "R": case(row) 8'b11110000,8'b10001000,8'b11110000,8'b10010000,8'b10001000,8'b10001000,8'b00000000,8'b00000000; endcase
            "O": case(row) 8'b01110000,8'b10001000,8'b10001000,8'b10001000,8'b10001000,8'b01110000,8'b00000000,8'b00000000; endcase
            "G": case(row) 8'b01110000,8'b10001000,8'b10000000,8'b10111000,8'b10001000,8'b01110000,8'b00000000,8'b00000000; endcase
            "A": case(row) 8'b01100000,8'b10010000,8'b10010000,8'b11110000,8'b10010000,8'b10010000,8'b00000000,8'b00000000; endcase
            "M": case(row) 8'b10001000,8'b11011000,8'b10101000,8'b10001000,8'b10001000,8'b10001000,8'b00000000,8'b00000000; endcase
            "C": case(row) 8'b01110000,8'b10001000,8'b10000000,8'b10000000,8'b10001000,8'b01110000,8'b00000000,8'b00000000; endcase
            "U": case(row) 8'b10001000,8'b10001000,8'b10001000,8'b10001000,8'b10001000,8'b01110000,8'b00000000,8'b00000000; endcase
            "N": case(row) 8'b10001000,8'b11001000,8'b10101000,8'b10011000,8'b10001000,8'b10001000,8'b00000000,8'b00000000; endcase
            "T": case(row) 8'b11111000,8'b00100000,8'b00100000,8'b00100000,8'b00100000,8'b00100000,8'b00000000,8'b00000000; endcase
            "E": case(row) 8'b11111000,8'b10000000,8'b11100000,8'b10000000,8'b10000000,8'b11111000,8'b00000000,8'b00000000; endcase
            " ": case(row) 8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000,8'b00000000; endcase
            default: pixels = 8'b00000000;
        endcase
    end
endmodule
